package pack;
import uvm_pkg::*;

`include "sequence_item.sv"
 `include "sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
endpackage
